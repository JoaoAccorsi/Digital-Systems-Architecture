// Structural Varilog implementation for expression Y = AB

module activity_2_structural_design (A, B, Y);

input A, B;
output Y;

and U1 (S, A, B);

endmodule
